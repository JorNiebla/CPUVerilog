module uc(input wire [15:0] opcode, input wire z, carry, output reg s_inc, s_inm, we3, wez, push, pop, output reg [2:0] op_alu);

  assign op_alu = opcode[26:24];
  assign s_inm = opcode[27];

  always @(opcode)
  begin
    s_inc = 1'b1;
    wez = 1'b0;
    we3 = 1'b0;
    push = 1'b0;
    pop = 1'b0;
    casez (opcode)
      16'b101?????????????: begin
        wez = z;
        we3 = 1'b1;
      end
      16'b100?????????????: begin
        we3 = 1'b1;
      end
      16'b11??????????????: begin
        we3 = 1'b1;
      end
      16'b01???????????01?: begin
        wez = z;
        we3 = 1'b1;
      end
      16'b01???????????00?: begin
        we3 = 1'b1;
      end
      16'b01???????????1??: begin
        we3 = 1'b1;
      end
      16'b001??????????000: begin //J
        s_inc = 1'b0;
      end
      16'b001??????????001: begin //JZ
        s_inc = ~z;
        
      end
      16'b001??????????010: begin //JNZ
        s_inc = z;
      end
      16'b001??????????011: begin //JA
        s_inc = ~z & ~carry;
      end
      16'b001??????????100: begin //JAE
        s_inc = carry;
      end
      16'b001??????????101: begin //JB
        s_inc = ~carry;
      end
      16'b001??????????110: begin //CALL
        s_inc = 1'b0;
        push = 1'b1;
      end
      16'b001??????????111: begin //RET
        pop = 1'b1;
      end
      16'b0001?????????011: begin //CMP
        wez = z;
      end
    endcase
  end

endmodule