module uc(input wire [5:0] opcode, input wire z, output reg s_inc, s_inm, we3, wez, push, pop, inm, carry, output reg [2:0] op_alu);

  initial begin
    we3 = 1'b0;

  end


endmodule